package svm_pkg;
    `include "svm_component.svh"
    `include "svm_factory.svh"
    `include "svm_registry.svh"
endpackage